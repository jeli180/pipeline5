//send hardcoded circle, line, square pixel data in software
//load weights based on mlp model outputs
//check if inference model worked by checking registers

