module dpu (
  input logic clk, rst,

  //from mmio
  input logic req, load,
  input logic [31:0] addr, write_data,

  //to mmio
  output logic ack, 
  output logic [31:0] read_data,

  //to screen
  output logic rd, wr, rs, cs, //rd, wr, cs are low active

  //from screen
  input logic interrupt, //low active

  inout wire [7:0] db
);

  /* RA8875 DPU description
      - mmio read/write cycle is when req goes high, load/addr/write_data are details of the
        transaction
      - every mmio transaction modeled as a dcache hit, so ack goes high the next cycle with 
        read_data if transaction is a read
      - using 8080 8b parrallel to interface with screen, all signals correspond to those in
        datasheet
      - db driven by both screen and this module, so modeled as wire
  */

  typedef enum {
    IDLE_C,
    INIT,
    CLEAR,
    POLL_INT,
    COORD,
    DRAW,
    SEND,
    WAIT_RECIEVE,
    WAIT_INFERENCE,
    PREP_CLEAR,
    FIX,
    DONE,
    CURSOR_RST,
    FULL_DONE
  } state_control;

  state_control stateC, next_stateC;

  typedef enum {
    IDLE_I,
    PREP_REG,
    PREP_REG2,
    INIT_REG,
    SEND_REG,
    END_REG,
    FINISH_REG,
    PREP_DATA,
    INIT_DATA,
    DATA,
    LAG_DATA,
    END_DATA,
    FINISH_DATA
  } state_interface;

  state_interface stateI, next_stateI;

  /* db is tri state
      - when i drive, i set drive high and set db_w
      - when drive is low, display is free to write to db, and i read db_r value
      - drive is default low;
  */

  logic [7:0] next_db_w, db_w;
  logic drive, next_drive, next_rs, next_cs, next_rd, next_wr;
  wire [7:0] db_r;

  assign db = drive ? db_w : 'z;
  assign db_r = db;

  //fsm control signals
  logic [18:0] ct, next_ct; //max ct number used is the total pixels (384,000)
  logic if_busy, next_if_busy;
  logic [7:0] screen_reg, screen_data, next_screen_reg, next_screen_data;
  logic screen_r, next_screen_r;
  logic [9:0] touchX, touchY, next_touchX, next_touchY, touchX3, touchY3; //stores touch coord to write to|technically Y doesn't need 10 bits
  //also using touchX, touchY as markers for active window origin during SEND to save space 
  logic [4:0] pixelbit, next_pixelbit; //tracks which bit of pixel_data we are on during SEND phase

  //register signals for outputs to CPU
  logic [31:0] next_shape, next_pixel_data, shape, pixel_data, full_done, next_full_done;
  logic [15:0] next_store, store; //store all shape data with valid bits
  logic next_ack;
  logic [31:0] next_read_data;

  //LINES CHANGED FOR SIM: 280, 428

  always_comb begin

    //mmio defaults
    next_ack = 0;
    next_read_data = '0; //next read data sent to cpu, synced with ack

    //registered values defaults
    next_shape = shape; //stores cpu sent shape data
    next_pixel_data = pixel_data; //generated by SEND state of control fsm
    next_full_done = full_done;

    //mmio req logic
    if (req) begin
      next_ack = 1;
      if (load) begin
        if (addr == 32'd4) next_read_data = pixel_data;
        else if (addr == 32'd8) next_read_data = full_done;
      end else begin
        if (addr == 32'd8) next_shape = write_data;
      end
    end

    //control fsm defaults
    next_ct = ct;
    next_if_busy = if_busy;
    next_screen_reg = screen_reg; //control fsm stores destination register to write/read to and from 
    next_screen_data = screen_data; //control fsm stores write data, interface fsm stores read data
    next_screen_r = screen_r; //control fsm stores whether to read/write to screen
    next_touchX = touchX; //registered x coord read from touch event by COORD state and used in DRAW state
    next_touchY = touchY;
    next_pixelbit = pixelbit;
    next_store = store;
    next_stateC = stateC;
    next_stateI = stateI;

    touchX3 = touchX + 10'd3;
    touchY3 = touchY + 10'd3;

    case (stateC) 
      IDLE_C: if (req && !load && addr == 32'd4) next_stateC = INIT; //transition on cpu signal
      INIT: begin
        if (!if_busy && stateI == IDLE_I) begin //double check, !if_busy should guarantee second condition
          if (ct > 18) begin //if ct is 19, initialization sequence is done
            next_stateC = CLEAR;
            next_ct = '0;
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;
            case (ct) //0-26 requests for interface fsm

              //sw reset
              19'd0: begin
                next_screen_reg = 8'h01;
                next_screen_data = 8'b00000001;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd1: begin
                next_screen_data = 8'b0;
                next_screen_r = 0;
                next_stateI = PREP_DATA;
              end

              //screen width and timing values
              19'd2: begin
                next_screen_reg = 8'h14;
                next_screen_data = 8'h63;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd3: begin
                next_screen_reg = 8'h16;
                next_screen_data = 8'h1F;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd4: begin
                next_screen_reg = 8'h17;
                next_screen_data = 8'h4;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd5: begin
                next_screen_reg = 8'h18;
                next_screen_data = 8'hF;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd6: begin
                next_screen_reg = 8'h19;
                next_screen_data = 8'hDF;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd7: begin
                next_screen_reg = 8'h1A;
                next_screen_data = 8'h1;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd8: begin
                next_screen_reg = 8'h1B;
                next_screen_data = 8'h2C;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd9: begin
                next_screen_reg = 8'h1D;
                next_screen_data = 8'h7;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd10: begin
                next_screen_reg = 8'h1F;
                next_screen_data = 8'h1;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end

              //turn display on
              19'd11: begin
                next_screen_reg = 8'h1;
                next_screen_data = 8'h80;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end

              //touchpad config
              19'd12: begin
                next_screen_reg = 8'h70;
                next_screen_data = 8'h80;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd13: begin
                next_screen_reg = 8'h71;
                next_screen_data = 8'h84;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end

              //interrupt enable
              19'd14: begin
                next_screen_reg = 8'hF0;
                next_screen_data = 8'h04;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end

              //set active window
              19'd15: begin
                next_screen_reg = 8'h34;
                next_screen_data = 8'h20;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd16: begin
                next_screen_reg = 8'h35;
                next_screen_data = 8'h03;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd17: begin
                next_screen_reg = 8'h36;
                next_screen_data = 8'hE0;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd18: begin
                next_screen_reg = 8'h37;
                next_screen_data = 8'h01;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              default:;
            endcase
          end
        end
      end
      CLEAR: begin
        if (!if_busy && stateI == IDLE_I) begin //double check, !if_busy should guarantee second condition
          //if (ct > 9) begin //simulation version
          if (ct > 383999) begin
            if (&store[15:12]) next_stateC = FIX;
            else next_stateC = POLL_INT;
            next_ct = '0;
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;

            if (ct == 0) begin
              next_screen_reg = 8'h2;
              next_screen_data = 8'b11111111;
              next_screen_r = 0;
              next_stateI = PREP_REG;
            end else begin
              next_stateI = PREP_DATA;
              //other values have stayed the same since ct = 0
            end
          end
        end
      end
      POLL_INT: if (!interrupt) next_stateC = COORD;
      COORD: begin
        //read from 72, 73, 74 to get coords, store the coords
        //if store high 4 bits on, shapes are already drawn, waiting for done signal from user
        if (!if_busy && stateI == IDLE_I) begin
          if (ct > 3) begin
            next_ct = '0;
            if (touchX > 480) begin
              if (&store[15:12]) next_stateC = CURSOR_RST;
              else next_stateC = SEND;
              next_touchX = '0;
              next_touchY = '0;
            end
            else begin
              if (&store[15:12]) next_stateC = POLL_INT;
              else next_stateC = DRAW;
            end
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;

            case (ct) 
              19'd0: begin
                next_screen_reg = 8'h72;
                next_screen_r = 1;
                next_stateI = PREP_REG;
              end
              19'd1: begin
                next_screen_reg = 8'h73;
                next_stateI = PREP_REG;
                //store the value interface FSM registered in screen_data before next transaction
                next_touchX = {screen_data, 2'b0};
              end
              19'd2: begin
                next_screen_reg = 8'h74;
                next_stateI = PREP_REG;
                next_touchY = {screen_data, 2'b0};
              end
              19'd3: begin //clear interrupt
                next_touchX = {touchX[9:2], screen_data[3:2]};
                next_touchY = {touchY[9:2], screen_data[1:0]};
                next_screen_reg = 8'hF1;
                next_screen_r = 0;
                next_stateI = PREP_REG;
                next_screen_data = 8'b00000100;
              end 
              default:;
            endcase
          end
        end
      end
      DRAW: begin
        //write mem cursor loc and stream black pixel to 2h
        if (!if_busy && stateI == IDLE_I) begin
          if (ct > 4) begin
            next_stateC = POLL_INT;
            next_ct = '0;
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;

            case (ct) 
              19'd0: begin
                next_screen_reg = 8'h46;
                next_screen_data = touchX[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd1: begin
                next_screen_reg = 8'h47;
                next_screen_data = {6'b0, touchX[9:8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd2: begin
                next_screen_reg = 8'h48;
                next_screen_data = touchY[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd3: begin
                next_screen_reg = 8'h49;
                next_screen_data = {7'b0, touchY[8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd4: begin
                next_screen_reg = 8'h2;
                next_screen_data = 8'b0;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              default:;
            endcase
          end
        end
      end
      SEND: begin
        /*
          - one bit of pixel_data is the product of ORing all pixels in a 4x4 block
          - pixel_data is filled with the 4x4 starting top left of each quadrant, 
            shifting to the right then down when finished with the row (similar to mem cursor)
        */
        if (!if_busy && stateI == IDLE_I) begin
          if (ct > 28) begin
            next_ct = '0;
            next_pixel_data[pixelbit] = pixel_data[pixelbit] || screen_data == 8'b0; //process last read data

            //check whether data bus is full
            if (pixelbit == 5'd29) begin
              next_pixelbit = '0;
              next_pixel_data[30] = 1'b1; //tells CPU data is valid
              next_stateC = WAIT_RECIEVE;
            end else begin
              next_pixelbit = pixelbit + 5'b1;
            end

            //need to keep at bottom for override
            if (touchX == 10'd236 && touchY == 10'd236) begin //first quad done
              next_touchX = 10'd240;
              next_touchY = '0;
            end else if (touchX == 10'd476 && touchY == 10'd236) begin //second quad done
              next_touchX = '0;
              next_touchY = 10'd240;
            end else if (touchX == 10'd236 && touchY == 10'd476) begin //third quad done
              next_touchX = 10'd240;
              next_touchY = 10'd240;
            end else if (touchX == 10'd476 && touchY == 10'd476) begin //all quads done, SEND state done
            //end else if (touchX == 10'd236 && touchY == 10'd12) begin //speed up simulation
              next_touchX = '0;
              next_touchY = '0;
              next_pixel_data[31] = 1'b1;
            end else if (touchX == 10'd236) begin
              next_touchX = '0;
              next_touchY = touchY + 4;
            end else if (touchX == 10'd476) begin
              next_touchX = 10'd240;
              next_touchY = touchY + 4;
            end else next_touchX = touchX + 4;

          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;

            case (ct)
              //0-7 to set active window according to pixelbit, touchX, touchY
              19'd0: begin
                next_screen_reg = 8'h30;
                next_screen_data = touchX[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end  
              19'd1: begin
                next_screen_reg = 8'h31;
                next_screen_data = {6'b0, touchX[9:8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd2: begin
                next_screen_reg = 8'h32;
                next_screen_data = touchY[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd3: begin
                next_screen_reg = 8'h33;
                next_screen_data = {7'b0, touchY[8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd4: begin
                next_screen_reg = 8'h34;
                next_screen_data = touchX3[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd5: begin
                next_screen_reg = 8'h35;
                next_screen_data = {6'b0, touchX3[9:8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd6: begin
                next_screen_reg = 8'h36;
                next_screen_data = touchY3[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd7: begin
                next_screen_reg = 8'h37;
                next_screen_data = {7'b0, touchY3[8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              //8-11 to set mem read cursor location
              19'd8: begin
                next_screen_reg = 8'h4A;
                next_screen_data = touchX[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd9: begin
                next_screen_reg = 8'h4B;
                next_screen_data = {6'b0, touchX[9:8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd10: begin
                next_screen_reg = 8'h4C;
                next_screen_data = touchY[7:0];
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd11: begin
                next_screen_reg = 8'h4D;
                next_screen_data = {7'b0, touchY[8]};
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end 
              //start sending pixels, d13 is different from default case as there is no data in screen_data
              //d12 because datasheet says there is a dummy read
              19'd12: begin
                next_screen_reg = 8'h2;
                next_screen_r = 1;
                next_stateI = PREP_REG;
              end
              19'd13: next_stateI = PREP_REG;
              default: begin
                next_stateI = PREP_DATA;
                //OR the bit of pixel_data with any bit of screen_data
                next_pixel_data[pixelbit] = pixel_data[pixelbit] || screen_data == 8'b0;
              end 
            endcase
          end
        end
      end
      WAIT_RECIEVE: begin
        if (req && !load && addr == 32'd4) begin
          next_pixel_data = '0;
          if (pixel_data[31]) next_stateC = WAIT_INFERENCE;
          else next_stateC = SEND;
        end
      end
      WAIT_INFERENCE: begin 
        //store all shape data in pixel bit, 4 msb are valids for each quadrant, 
        //transition when all 4msb are high
        if (&store[15:12]) next_stateC = PREP_CLEAR;
        case (shape[6:3])
          4'b0001: begin 
            next_store[12] = 1'b1;
            next_store[2:0] = shape[2:0];
          end
          4'b0010: begin
            next_store[13] = 1'b1;
            next_store[5:3] = shape[2:0];
          end
          4'b0100: begin
            next_store[14] = 1'b1;
            next_store[8:6] = shape[2:0];
          end
          4'b1000: begin
            next_store[15] = 1'b1;
            next_store[11:9] = shape[2:0];
          end
          default:;
        endcase
      end
      PREP_CLEAR: begin
        if (!if_busy && stateI == IDLE_I) begin
          if (ct > 7) begin 
            next_stateC = CLEAR;
            next_ct = '0;
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;

            case (ct)
              //0-7 set active window
              19'd0: begin
                next_screen_reg = 8'h30;
                next_screen_data = 8'b0;
                next_screen_r = 0;
                next_stateI = PREP_REG;
              end
              19'd1: begin
                next_screen_reg = 8'h31;
                next_screen_data = 8'b0;
                next_stateI = PREP_REG;
              end
              19'd2: begin
                next_screen_reg = 8'h32;
                next_screen_data = 8'b0;
                next_stateI = PREP_REG;
              end
              19'd3: begin
                next_screen_reg = 8'h33;
                next_screen_data = 8'b0;
                next_stateI = PREP_REG;
              end
              19'd4: begin
                next_screen_reg = 8'h34;
                next_screen_data = 8'b00100000;;
                next_stateI = PREP_REG;
              end
              19'd5: begin
                next_screen_reg = 8'h35;
                next_screen_data = 8'b00000011;
                next_stateI = PREP_REG;
              end
              19'd6: begin
                next_screen_reg = 8'h36;
                next_screen_data = 8'b01110000;
                next_stateI = PREP_REG;
              end
              19'd7: begin
                next_screen_reg = 8'h37;
                next_screen_data = 8'b1;
                next_stateI = PREP_REG;
              end
              default:;
            endcase
          end
        end
      end  
      FIX: begin //100 is circle, 010 is square, 001 is line
        if (!if_busy && stateI == IDLE_I) begin
          if (ct > 8) begin 
            next_stateC = DONE;
            next_ct = '0;
            next_screen_data = 8'b1100000; //significant to DONE state
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;

            case (ct) 
              //use 45h as a dummy reg to write to

              //circle center and line/square horizontal start coord
              19'd0: begin
                next_screen_r = 0;
                next_stateI = PREP_REG;
                if (store[12]) begin
                  next_screen_data = store[2] ? 8'b01110111 : 8'b00111011;
                  next_screen_reg = store[2] ? 8'h99 : 8'h91;
                end else if (store[13]) begin 
                  next_screen_data = store[5] ? 8'b01100111 : 8'b00101011;
                  next_screen_reg = store[5] ? 8'h99 : 8'h91;
                end else if (store[14]) begin 
                  next_screen_data = store[8] ? 8'b01110111 : 8'b00111011;
                  next_screen_reg = store[8] ? 8'h99 : 8'h91;
                end else if (store[15]) begin 
                  next_screen_data = store[11] ? 8'b01100111 : 8'b00101011;
                  next_screen_reg = store[11] ? 8'h99 : 8'h91;
                end
              end
              19'd1: begin
                next_stateI = PREP_REG;
                if (store[12]) begin 
                  next_screen_data = 8'b0;
                  next_screen_reg = store[2] ? 8'h9A : 8'h92;
                end else if (store[13]) begin
                  next_screen_data = 8'b1;
                  next_screen_reg = store[5] ? 8'h9A : 8'h92;
                end else if (store[14]) begin
                  next_screen_data = 8'b0;
                  next_screen_reg = store[8] ? 8'h9A : 8'h92;
                end else if (store[15]) begin
                  next_screen_data = 8'b1;
                  next_screen_reg = store[11] ? 8'h9A : 8'h92;
                end
              end

              //circle center and line/square vertical start coord
              19'd2: begin
                next_stateI = PREP_REG;
                if (store[12]) begin
                  next_screen_data = store[2] ? 8'b01110111 : 8'b00111011;
                  next_screen_reg = store[2] ? 8'h9B : 8'h93;
                end else if (store[13]) begin 
                  next_screen_data = store[5] ? 8'b01110111 : 8'b00111011;
                  next_screen_reg = store[2] ? 8'h9B : 8'h93;
                end else if (store[14]) begin
                  next_screen_data = store[8] ? 8'b01100111 : 8'b00101011;
                  next_screen_reg = store[8] ? 8'h9B : 8'h93;
                end else if (store[15]) begin
                  next_screen_data = store[11] ? 8'b01100111 : 8'b00101011;
                  next_screen_reg = store[11] ? 8'h9B : 8'h93;
                end
              end 
              19'd3: begin
                next_stateI = PREP_REG;
                if (store[12]) begin 
                  next_screen_data = 8'b0;
                  next_screen_reg = store[2] ? 8'h9C : 8'h94;
                end else if (store[13]) begin
                  next_screen_data = 8'b0;
                  next_screen_reg = store[5] ? 8'h9C : 8'h94;
                end else if (store[14]) begin
                  next_screen_data = 8'b1;
                  next_screen_reg = store[8] ? 8'h9C : 8'h94;
                end else if (store[15]) begin
                  next_screen_data = 8'b1;
                  next_screen_reg = store[11] ? 8'h9C : 8'h94;
                end
              end

              //circle radius for first only, square/line horizontal end coord
              19'd4: begin
                next_stateI = PREP_REG;
                if (store[12]) begin
                  next_screen_data = store[2] ? 8'b01010000 : 8'b10110011;
                  next_screen_reg = store[2] ? 8'h9D : 8'h95;
                end else if (store[13]) begin
                  next_screen_data = store[5] ? 8'b01010000 : 8'b10100011;
                  next_screen_reg = store[5] ? 8'h9D : 8'h95;
                end else if (store[14]) begin
                  next_screen_data = store[8] ? 8'b01010000 : 8'b10110011;
                  next_screen_reg = store[8] ? 8'h9D : 8'h95;
                end else if (store[15]) begin
                  next_screen_data = store[11] ? 8'b01010000 : 8'b10100011;
                  next_screen_reg = store[11] ? 8'h9D : 8'h95;
                end
              end
              19'd5: begin
                next_stateI = PREP_REG;
                if (store[12]) begin
                  next_screen_data = 8'b0;
                  next_screen_reg = store[2] ? 8'h45 : 8'h96;
                end else if (store[13]) begin
                  next_screen_data = store[5] ? 8'b0 : 8'b1;
                  next_screen_reg = store[5] ? 8'h45 : 8'h96;
                end else if (store[14]) begin
                  next_screen_data = 8'b0;
                  next_screen_reg = store[8] ? 8'h45 : 8'h96;
                end else if (store[15]) begin
                  next_screen_data = store[11] ? 8'b0 : 8'b1;
                  next_screen_reg = store[11] ? 8'h45 : 8'h96;
                end
              end

              //square/line vertical end coord
              19'd6: begin
                next_stateI = PREP_REG;
                if (store[12]) begin
                  next_screen_data = store[2] ? 8'b0 : 8'b10110011;
                  next_screen_reg = store[2] ? 8'h45 : 8'h97;
                end else if (store[13]) begin
                  next_screen_data = store[5] ? 8'b0 : 8'b10110011;
                  next_screen_reg = store[5] ? 8'h45 : 8'h97;
                end else if (store[14]) begin
                  next_screen_data = store[8] ? 8'b0 : 8'b10100011;
                  next_screen_reg = store[8] ? 8'h45 : 8'h97;
                end else if (store[15]) begin
                  next_screen_data = store[11] ? 8'b0 : 8'b10100011;
                  next_screen_reg = store[11] ? 8'h45 : 8'h97;
                end
              end
              19'd7: begin
                next_stateI = PREP_REG;
                if (store[12]) begin 
                  next_screen_data = 8'b0;
                  next_screen_reg = store[2] ? 8'h45 : 8'h98;
                end else if (store[13]) begin
                  next_screen_data = 8'b0;
                  next_screen_reg = store[5] ? 8'h45 : 8'h98;
                end else if (store[14]) begin
                  next_screen_data = store[8] ? 8'b0 : 8'b1;
                  next_screen_reg = store[8] ? 8'h45 : 8'h98;
                end else if (store[15]) begin
                  next_screen_data = store[11] ? 8'b0 : 8'b1;
                  next_screen_reg = store[11] ? 8'h45 : 8'h98;
                end
              end

              //start draw reg
              19'd8: begin
                next_screen_reg = 8'h90;
                next_stateI = PREP_REG;
                if (store[12]) begin
                  next_screen_data = store[2] ? 8'b01000000 : 
                                     store[1] ? 8'b10010000 : //square
                                                8'b10000000 ;
                end else if (store[13]) begin
                  next_screen_data = store[5] ? 8'b01000000 : 
                                     store[4] ? 8'b10010000 : 
                                                8'b10000000 ;
                end else if (store[14]) begin
                  next_screen_data = store[8] ? 8'b01000000 : 
                                     store[7] ? 8'b10010000 : 
                                                8'b10000000 ;
                end else if (store[15]) begin
                  next_screen_data = store[11] ? 8'b01000000 : 
                                     store[10] ? 8'b10010000 : 
                                                 8'b10000000 ;
                end
              end
              default:;
            endcase
          end
        end
      end
      DONE: begin
        //update store after each shape done printing
        //transition to CURSOR_RST when all shapes done printing
        if (!if_busy && stateI == IDLE_I) begin 
          if (!screen_data[7] && !screen_data[6]) begin //checks if draw function done
            if (store[12]) begin
              next_store = {4'b1110, store[11:3], 3'b0};
              next_stateC = FIX;
            end else if (store[13]) begin
              next_store = {4'b1100, store[11:6], 6'b0};
              next_stateC = FIX;
            end else if (store[14]) begin
              next_store = {4'b1000, store[11:9], 9'b0};
              next_stateC = FIX;
            end else begin
              next_store = 16'hF000; //set up correct COORD state behavior
              next_stateC = POLL_INT; //POLL_INT waits for user to clear shapes
            end
          end else begin
            next_if_busy = 1;
            next_stateI = PREP_REG;
            next_screen_reg = 8'h90;
            next_screen_r = 1'b1;
          end
        end
      end
      CURSOR_RST: begin
        //reset all tracking registers: pixel_data, ct, screen_data, screen_reg, screen_r,
        //touchX, touchY, pixelbit 
        //reset mem cursor location, read is automatically set within the statemachine to default
        //46-49
        if (!if_busy && stateI == IDLE_I) begin 
          if (ct > 3) begin 
            next_stateC = FULL_DONE;
            next_ct = '0;
            next_pixel_data = '0;
            next_screen_data = '0;
            next_screen_reg = '0;
            next_touchX = '0;
            next_touchY = '0;
            next_pixelbit = '0;
            next_store = '0;
          end else begin
            next_ct = ct + 19'b1;
            next_if_busy = 1;
            next_screen_data = '0;

            //reset mem write cursor
            case (ct) 
              19'd0: begin
                next_screen_reg = 8'h46;
                next_screen_r = 1'b0;
                next_stateI = PREP_REG;
              end
              19'd1: begin
                next_screen_reg = 8'h47;
                next_stateI = PREP_REG;
              end
              19'd2: begin
                next_screen_reg = 8'h48;
                next_stateI = PREP_REG;
              end
              19'd3: begin
                next_screen_reg = 8'h49;
                next_stateI = PREP_REG;
              end
              default:;
            endcase
          end
        end
      end
      FULL_DONE: begin //fill full done register that CPU polls by loading from h8, cpu acks by h4 store
        next_full_done = 32'd1;
        if (req && !load && addr == 32'd4) begin
          next_stateC = CLEAR;
          next_full_done = '0;
        end
      end
      default:;
    endcase
    
    //interface signal defaults
    next_rd = 1;
    next_wr = 1;
    next_rs = 1;
    next_cs = 1;
    next_drive = 0;
    next_db_w = '0;

    case (stateI)
      PREP_REG: begin
        next_stateI = PREP_REG2;
      end
      PREP_REG2: begin
        next_cs = 0;
        next_stateI = INIT_REG;
      end
      INIT_REG: begin
        next_cs = 0;
        next_wr = 0;
        next_stateI = SEND_REG;
      end
      SEND_REG: begin
        next_cs = 0;
        next_wr = 0;
        next_drive = 1;
        next_db_w = screen_reg;
        next_stateI = END_REG;
      end
      END_REG: begin
        next_cs = 0;
        next_stateI = FINISH_REG;
      end
      FINISH_REG: begin
        next_rs = 0;
        next_stateI = PREP_DATA;
      end
      PREP_DATA: begin
        next_cs = 0;
        next_rs = 0;
        next_stateI = INIT_DATA;
      end
      INIT_DATA: begin
        next_cs = 0;
        next_rs = 0;
        if (screen_r) next_rd = 0;
        else next_wr = 0;
        next_stateI = DATA;
      end
      DATA: begin
        next_cs = 0;
        next_rs = 0;
        if (screen_r) begin
          next_rd = 0;
        end else begin
          next_wr = 0;
          next_drive = 1;
          next_db_w = screen_data;
        end
        next_stateI = LAG_DATA;
      end
      LAG_DATA: begin
        next_cs = 0;
        next_rs = 0;
        if (screen_r) begin
          next_rd = 0;
          next_screen_data = db_r;
        end else begin
          next_wr = 0;
          next_drive = 1;
          next_db_w = screen_data;
        end
        next_stateI = END_DATA;
      end
      END_DATA: begin
        next_cs = 0;
        next_rs = 0;
        next_stateI = FINISH_DATA;
      end
      FINISH_DATA: begin
        next_if_busy = 0;
        next_stateI = IDLE_I;
      end
      default:;
    endcase
  end 

  always_ff @(posedge clk, posedge rst) begin
    if (rst) begin
      ct <= '0;
      if_busy <= 0;
      screen_reg <= '0;
      screen_data <= '0;
      screen_r <= 0;
      touchX <= '0;
      touchY <= '0;
      pixelbit <= '0;
      shape <= '0;
      pixel_data <= '0;
      store <= '0;
      ack <= 0;
      read_data <= '0;
      cs <= 1'b1;
      rs <= 1'b1;
      wr <= 1'b1;
      rd <= 1'b1;
      drive <= 0;
      db_w <= '0;
      full_done <= '0;
      stateC <= IDLE_C;
      stateI <= IDLE_I;
    end else begin
      ct <= next_ct;
      if_busy <= next_if_busy;
      screen_reg <= next_screen_reg;
      screen_data <= next_screen_data;
      screen_r <= next_screen_r;
      touchX <= next_touchX;
      touchY <= next_touchY;
      pixelbit <= next_pixelbit;
      shape <= next_shape;
      pixel_data <= next_pixel_data;
      store <= next_store;
      ack <= next_ack;
      read_data <= next_read_data;
      cs <= next_cs;
      rs <= next_rs;
      wr <= next_wr;
      rd <= next_rd;
      drive <= next_drive;
      db_w <= next_db_w;
      full_done <= next_full_done;
      stateC <= next_stateC;
      stateI <= next_stateI;
    end
  end

endmodule